code,name,start_date,end_date,days,p_change
603118,共进股份,2019-10-25,2019-10-18,5,0
002815,崇达技术,2019-11-08,2019-11-01,5,0
002756,永兴材料,2019-11-08,2019-11-01,5,0
603386,广东骏亚,2019-11-08,2019-11-01,5,0
603133,碳元科技,2019-11-08,2019-11-01,5,0
603799,华友钴业,2019-11-08,2019-11-01,5,0
002587,奥拓电子,2019-10-25,2019-10-18,5,0
603060,国检集团,2019-11-08,2019-11-01,5,0
603920,世运电路,2019-11-01,2019-10-25,5,0
002855,捷荣技术,2019-11-08,2019-11-01,5,0
600845,宝信软件,2019-11-08,2019-11-01,5,0
600882,妙可蓝多,2019-11-08,2019-11-01,5,0
002683,宏大爆破,2019-10-25,2019-10-18,5,0
002185,华天科技,2019-11-01,2019-10-25,5,0
000673,当代东方,2019-11-08,2019-11-01,5,0
603881,数据港,2019-11-08,2019-11-01,5,0
002138,顺络电子,2019-11-08,2019-11-01,5,0
603228,景旺电子,2019-11-08,2019-11-01,5,0
002808,恒久科技,2019-11-01,2019-10-25,5,0
603136,天目湖,2019-10-18,2019-10-11,5,0
603180,金牌厨柜,2019-11-01,2019-10-25,5,0
600818,中路股份,2019-10-25,2019-10-18,5,0
000977,浪潮信息,2019-10-25,2019-10-18,5,0
002129,中环股份,2019-11-08,2019-11-01,5,0
600093,易见股份,2019-10-25,2019-10-18,5,0
002414,高德红外,2019-11-08,2019-11-01,5,0
002528,英飞拓,2019-10-11,2019-09-30,5,0
002531,天顺风能,2019-11-08,2019-11-01,5,0
